module FontROM (
    input wire [7:0] char_code,
    input wire [2:0] row,
    output reg [7:0] pixels
);

    always @(*) begin
        case ({char_code, row})
            {8'd65, 3'd0}: pixels = 8'b00011000;
            {8'd65, 3'd1}: pixels = 8'b00100100;
            {8'd65, 3'd2}: pixels = 8'b01000010;
            {8'd65, 3'd3}: pixels = 8'b01111110;
            {8'd65, 3'd4}: pixels = 8'b01000010;
            {8'd65, 3'd5}: pixels = 8'b01000010;
            {8'd65, 3'd6}: pixels = 8'b01000010;
            {8'd65, 3'd7}: pixels = 8'b00000000;
            {8'd66, 3'd0}: pixels = 8'b01111100;
            {8'd66, 3'd1}: pixels = 8'b01000010;
            {8'd66, 3'd2}: pixels = 8'b01000010;
            {8'd66, 3'd3}: pixels = 8'b01111100;
            {8'd66, 3'd4}: pixels = 8'b01000010;
            {8'd66, 3'd5}: pixels = 8'b01000010;
            {8'd66, 3'd6}: pixels = 8'b01111100;
            {8'd66, 3'd7}: pixels = 8'b00000000;
            {8'd67, 3'd0}: pixels = 8'b00111100;
            {8'd67, 3'd1}: pixels = 8'b01000010;
            {8'd67, 3'd2}: pixels = 8'b01000000;
            {8'd67, 3'd3}: pixels = 8'b01000000;
            {8'd67, 3'd4}: pixels = 8'b01000000;
            {8'd67, 3'd5}: pixels = 8'b01000010;
            {8'd67, 3'd6}: pixels = 8'b00111100;
            {8'd67, 3'd7}: pixels = 8'b00000000;
            {8'd68, 3'd0}: pixels = 8'b01111000;
            {8'd68, 3'd1}: pixels = 8'b01000100;
            {8'd68, 3'd2}: pixels = 8'b01000010;
            {8'd68, 3'd3}: pixels = 8'b01000010;
            {8'd68, 3'd4}: pixels = 8'b01000010;
            {8'd68, 3'd5}: pixels = 8'b01000100;
            {8'd68, 3'd6}: pixels = 8'b01111000;
            {8'd68, 3'd7}: pixels = 8'b00000000;
            {8'd69, 3'd0}: pixels = 8'b01111110;
            {8'd69, 3'd1}: pixels = 8'b01000000;
            {8'd69, 3'd2}: pixels = 8'b01000000;
            {8'd69, 3'd3}: pixels = 8'b01111100;
            {8'd69, 3'd4}: pixels = 8'b01000000;
            {8'd69, 3'd5}: pixels = 8'b01000000;
            {8'd69, 3'd6}: pixels = 8'b01111110;
            {8'd69, 3'd7}: pixels = 8'b00000000;
            {8'd70, 3'd0}: pixels = 8'b01111110;
            {8'd70, 3'd1}: pixels = 8'b01000000;
            {8'd70, 3'd2}: pixels = 8'b01000000;
            {8'd70, 3'd3}: pixels = 8'b01111100;
            {8'd70, 3'd4}: pixels = 8'b01000000;
            {8'd70, 3'd5}: pixels = 8'b01000000;
            {8'd70, 3'd6}: pixels = 8'b01000000;
            {8'd70, 3'd7}: pixels = 8'b00000000;
            {8'd71, 3'd0}: pixels = 8'b00111100;
            {8'd71, 3'd1}: pixels = 8'b01000010;
            {8'd71, 3'd2}: pixels = 8'b01000000;
            {8'd71, 3'd3}: pixels = 8'b01001110;
            {8'd71, 3'd4}: pixels = 8'b01000010;
            {8'd71, 3'd5}: pixels = 8'b01000010;
            {8'd71, 3'd6}: pixels = 8'b00111100;
            {8'd71, 3'd7}: pixels = 8'b00000000;
            {8'd72, 3'd0}: pixels = 8'b01000010;
            {8'd72, 3'd1}: pixels = 8'b01000010;
            {8'd72, 3'd2}: pixels = 8'b01000010;
            {8'd72, 3'd3}: pixels = 8'b01111110;
            {8'd72, 3'd4}: pixels = 8'b01000010;
            {8'd72, 3'd5}: pixels = 8'b01000010;
            {8'd72, 3'd6}: pixels = 8'b01000010;
            {8'd72, 3'd7}: pixels = 8'b00000000;
            {8'd73, 3'd0}: pixels = 8'b00111100;
            {8'd73, 3'd1}: pixels = 8'b00001000;
            {8'd73, 3'd2}: pixels = 8'b00001000;
            {8'd73, 3'd3}: pixels = 8'b00001000;
            {8'd73, 3'd4}: pixels = 8'b00001000;
            {8'd73, 3'd5}: pixels = 8'b00001000;
            {8'd73, 3'd6}: pixels = 8'b00111100;
            {8'd73, 3'd7}: pixels = 8'b00000000;
            {8'd74, 3'd0}: pixels = 8'b00011110;
            {8'd74, 3'd1}: pixels = 8'b00000100;
            {8'd74, 3'd2}: pixels = 8'b00000100;
            {8'd74, 3'd3}: pixels = 8'b00000100;
            {8'd74, 3'd4}: pixels = 8'b01000100;
            {8'd74, 3'd5}: pixels = 8'b01000100;
            {8'd74, 3'd6}: pixels = 8'b00111000;
            {8'd74, 3'd7}: pixels = 8'b00000000;
            {8'd75, 3'd0}: pixels = 8'b01000010;
            {8'd75, 3'd1}: pixels = 8'b01000100;
            {8'd75, 3'd2}: pixels = 8'b01001000;
            {8'd75, 3'd3}: pixels = 8'b01110000;
            {8'd75, 3'd4}: pixels = 8'b01001000;
            {8'd75, 3'd5}: pixels = 8'b01000100;
            {8'd75, 3'd6}: pixels = 8'b01000010;
            {8'd75, 3'd7}: pixels = 8'b00000000;
            {8'd76, 3'd0}: pixels = 8'b01000000;
            {8'd76, 3'd1}: pixels = 8'b01000000;
            {8'd76, 3'd2}: pixels = 8'b01000000;
            {8'd76, 3'd3}: pixels = 8'b01000000;
            {8'd76, 3'd4}: pixels = 8'b01000000;
            {8'd76, 3'd5}: pixels = 8'b01000000;
            {8'd76, 3'd6}: pixels = 8'b01111110;
            {8'd76, 3'd7}: pixels = 8'b00000000;
            {8'd77, 3'd0}: pixels = 8'b01000010;
            {8'd77, 3'd1}: pixels = 8'b01100110;
            {8'd77, 3'd2}: pixels = 8'b01011010;
            {8'd77, 3'd3}: pixels = 8'b01011010;
            {8'd77, 3'd4}: pixels = 8'b01000010;
            {8'd77, 3'd5}: pixels = 8'b01000010;
            {8'd77, 3'd6}: pixels = 8'b01000010;
            {8'd77, 3'd7}: pixels = 8'b00000000;
            {8'd78, 3'd0}: pixels = 8'b01000010;
            {8'd78, 3'd1}: pixels = 8'b01100010;
            {8'd78, 3'd2}: pixels = 8'b01010010;
            {8'd78, 3'd3}: pixels = 8'b01001010;
            {8'd78, 3'd4}: pixels = 8'b01000110;
            {8'd78, 3'd5}: pixels = 8'b01000010;
            {8'd78, 3'd6}: pixels = 8'b01000010;
            {8'd78, 3'd7}: pixels = 8'b00000000;
            {8'd79, 3'd0}: pixels = 8'b00111100;
            {8'd79, 3'd1}: pixels = 8'b01000010;
            {8'd79, 3'd2}: pixels = 8'b01000010;
            {8'd79, 3'd3}: pixels = 8'b01000010;
            {8'd79, 3'd4}: pixels = 8'b01000010;
            {8'd79, 3'd5}: pixels = 8'b01000010;
            {8'd79, 3'd6}: pixels = 8'b00111100;
            {8'd79, 3'd7}: pixels = 8'b00000000;
            {8'd80, 3'd0}: pixels = 8'b01111100;
            {8'd80, 3'd1}: pixels = 8'b01000010;
            {8'd80, 3'd2}: pixels = 8'b01000010;
            {8'd80, 3'd3}: pixels = 8'b01111100;
            {8'd80, 3'd4}: pixels = 8'b01000000;
            {8'd80, 3'd5}: pixels = 8'b01000000;
            {8'd80, 3'd6}: pixels = 8'b01000000;
            {8'd80, 3'd7}: pixels = 8'b00000000;
            {8'd81, 3'd0}: pixels = 8'b00111100;
            {8'd81, 3'd1}: pixels = 8'b01000010;
            {8'd81, 3'd2}: pixels = 8'b01000010;
            {8'd81, 3'd3}: pixels = 8'b01000010;
            {8'd81, 3'd4}: pixels = 8'b01001010;
            {8'd81, 3'd5}: pixels = 8'b01000100;
            {8'd81, 3'd6}: pixels = 8'b00111010;
            {8'd81, 3'd7}: pixels = 8'b00000000;
            {8'd82, 3'd0}: pixels = 8'b01111100;
            {8'd82, 3'd1}: pixels = 8'b01000010;
            {8'd82, 3'd2}: pixels = 8'b01000010;
            {8'd82, 3'd3}: pixels = 8'b01111100;
            {8'd82, 3'd4}: pixels = 8'b01001000;
            {8'd82, 3'd5}: pixels = 8'b01000100;
            {8'd82, 3'd6}: pixels = 8'b01000010;
            {8'd82, 3'd7}: pixels = 8'b00000000;
            {8'd83, 3'd0}: pixels = 8'b00111100;
            {8'd83, 3'd1}: pixels = 8'b01000010;
            {8'd83, 3'd2}: pixels = 8'b01000000;
            {8'd83, 3'd3}: pixels = 8'b00111100;
            {8'd83, 3'd4}: pixels = 8'b00000010;
            {8'd83, 3'd5}: pixels = 8'b01000010;
            {8'd83, 3'd6}: pixels = 8'b00111100;
            {8'd83, 3'd7}: pixels = 8'b00000000;
            {8'd84, 3'd0}: pixels = 8'b01111111;
            {8'd84, 3'd1}: pixels = 8'b01001001;
            {8'd84, 3'd2}: pixels = 8'b00001000;
            {8'd84, 3'd3}: pixels = 8'b00001000;
            {8'd84, 3'd4}: pixels = 8'b00001000;
            {8'd84, 3'd5}: pixels = 8'b00001000;
            {8'd84, 3'd6}: pixels = 8'b00011100;
            {8'd84, 3'd7}: pixels = 8'b00000000;
            {8'd85, 3'd0}: pixels = 8'b01000010;
            {8'd85, 3'd1}: pixels = 8'b01000010;
            {8'd85, 3'd2}: pixels = 8'b01000010;
            {8'd85, 3'd3}: pixels = 8'b01000010;
            {8'd85, 3'd4}: pixels = 8'b01000010;
            {8'd85, 3'd5}: pixels = 8'b01000010;
            {8'd85, 3'd6}: pixels = 8'b00111100;
            {8'd85, 3'd7}: pixels = 8'b00000000;
            {8'd86, 3'd0}: pixels = 8'b01000010;
            {8'd86, 3'd1}: pixels = 8'b01000010;
            {8'd86, 3'd2}: pixels = 8'b01000010;
            {8'd86, 3'd3}: pixels = 8'b01000010;
            {8'd86, 3'd4}: pixels = 8'b00100100;
            {8'd86, 3'd5}: pixels = 8'b00100100;
            {8'd86, 3'd6}: pixels = 8'b00011000;
            {8'd86, 3'd7}: pixels = 8'b00000000;
            {8'd87, 3'd0}: pixels = 8'b01000010;
            {8'd87, 3'd1}: pixels = 8'b01000010;
            {8'd87, 3'd2}: pixels = 8'b01000010;
            {8'd87, 3'd3}: pixels = 8'b01011010;
            {8'd87, 3'd4}: pixels = 8'b01011010;
            {8'd87, 3'd5}: pixels = 8'b01100110;
            {8'd87, 3'd6}: pixels = 8'b01000010;
            {8'd87, 3'd7}: pixels = 8'b00000000;
            {8'd88, 3'd0}: pixels = 8'b01000010;
            {8'd88, 3'd1}: pixels = 8'b00100100;
            {8'd88, 3'd2}: pixels = 8'b00011000;
            {8'd88, 3'd3}: pixels = 8'b00011000;
            {8'd88, 3'd4}: pixels = 8'b00011000;
            {8'd88, 3'd5}: pixels = 8'b00100100;
            {8'd88, 3'd6}: pixels = 8'b01000010;
            {8'd88, 3'd7}: pixels = 8'b00000000;
            {8'd89, 3'd0}: pixels = 8'b01000010;
            {8'd89, 3'd1}: pixels = 8'b01000010;
            {8'd89, 3'd2}: pixels = 8'b00100100;
            {8'd89, 3'd3}: pixels = 8'b00011000;
            {8'd89, 3'd4}: pixels = 8'b00001000;
            {8'd89, 3'd5}: pixels = 8'b00001000;
            {8'd89, 3'd6}: pixels = 8'b00011100;
            {8'd89, 3'd7}: pixels = 8'b00000000;
            {8'd90, 3'd0}: pixels = 8'b01111110;
            {8'd90, 3'd1}: pixels = 8'b00000010;
            {8'd90, 3'd2}: pixels = 8'b00000100;
            {8'd90, 3'd3}: pixels = 8'b00001000;
            {8'd90, 3'd4}: pixels = 8'b00010000;
            {8'd90, 3'd5}: pixels = 8'b00100000;
            {8'd90, 3'd6}: pixels = 8'b01111110;
            {8'd90, 3'd7}: pixels = 8'b00000000;
            {8'd48, 3'd0}: pixels = 8'b00111100;
            {8'd48, 3'd1}: pixels = 8'b01100110;
            {8'd48, 3'd2}: pixels = 8'b01101110;
            {8'd48, 3'd3}: pixels = 8'b01110110;
            {8'd48, 3'd4}: pixels = 8'b01100110;
            {8'd48, 3'd5}: pixels = 8'b01100110;
            {8'd48, 3'd6}: pixels = 8'b00111100;
            {8'd48, 3'd7}: pixels = 8'b00000000;
            {8'd49, 3'd0}: pixels = 8'b00011000;
            {8'd49, 3'd1}: pixels = 8'b00111000;
            {8'd49, 3'd2}: pixels = 8'b00011000;
            {8'd49, 3'd3}: pixels = 8'b00011000;
            {8'd49, 3'd4}: pixels = 8'b00011000;
            {8'd49, 3'd5}: pixels = 8'b00011000;
            {8'd49, 3'd6}: pixels = 8'b00111100;
            {8'd49, 3'd7}: pixels = 8'b00000000;
            {8'd50, 3'd0}: pixels = 8'b00111100;
            {8'd50, 3'd1}: pixels = 8'b01100110;
            {8'd50, 3'd2}: pixels = 8'b00000110;
            {8'd50, 3'd3}: pixels = 8'b00001100;
            {8'd50, 3'd4}: pixels = 8'b00011000;
            {8'd50, 3'd5}: pixels = 8'b00110000;
            {8'd50, 3'd6}: pixels = 8'b01111110;
            {8'd50, 3'd7}: pixels = 8'b00000000;
            {8'd51, 3'd0}: pixels = 8'b00111100;
            {8'd51, 3'd1}: pixels = 8'b01100110;
            {8'd51, 3'd2}: pixels = 8'b00000110;
            {8'd51, 3'd3}: pixels = 8'b00011100;
            {8'd51, 3'd4}: pixels = 8'b00000110;
            {8'd51, 3'd5}: pixels = 8'b01100110;
            {8'd51, 3'd6}: pixels = 8'b00111100;
            {8'd51, 3'd7}: pixels = 8'b00000000;
            {8'd52, 3'd0}: pixels = 8'b00001100;
            {8'd52, 3'd1}: pixels = 8'b00011100;
            {8'd52, 3'd2}: pixels = 8'b00101100;
            {8'd52, 3'd3}: pixels = 8'b01001100;
            {8'd52, 3'd4}: pixels = 8'b01111110;
            {8'd52, 3'd5}: pixels = 8'b00001100;
            {8'd52, 3'd6}: pixels = 8'b00001100;
            {8'd52, 3'd7}: pixels = 8'b00000000;
            {8'd53, 3'd0}: pixels = 8'b01111110;
            {8'd53, 3'd1}: pixels = 8'b01100000;
            {8'd53, 3'd2}: pixels = 8'b01111100;
            {8'd53, 3'd3}: pixels = 8'b00000110;
            {8'd53, 3'd4}: pixels = 8'b00000110;
            {8'd53, 3'd5}: pixels = 8'b01100110;
            {8'd53, 3'd6}: pixels = 8'b00111100;
            {8'd53, 3'd7}: pixels = 8'b00000000;
            {8'd54, 3'd0}: pixels = 8'b00011100;
            {8'd54, 3'd1}: pixels = 8'b00110000;
            {8'd54, 3'd2}: pixels = 8'b01100000;
            {8'd54, 3'd3}: pixels = 8'b01111100;
            {8'd54, 3'd4}: pixels = 8'b01100110;
            {8'd54, 3'd5}: pixels = 8'b01100110;
            {8'd54, 3'd6}: pixels = 8'b00111100;
            {8'd54, 3'd7}: pixels = 8'b00000000;
            {8'd55, 3'd0}: pixels = 8'b01111110;
            {8'd55, 3'd1}: pixels = 8'b00000110;
            {8'd55, 3'd2}: pixels = 8'b00001100;
            {8'd55, 3'd3}: pixels = 8'b00011000;
            {8'd55, 3'd4}: pixels = 8'b00110000;
            {8'd55, 3'd5}: pixels = 8'b00110000;
            {8'd55, 3'd6}: pixels = 8'b00110000;
            {8'd55, 3'd7}: pixels = 8'b00000000;
            {8'd56, 3'd0}: pixels = 8'b00111100;
            {8'd56, 3'd1}: pixels = 8'b01100110;
            {8'd56, 3'd2}: pixels = 8'b01100110;
            {8'd56, 3'd3}: pixels = 8'b00111100;
            {8'd56, 3'd4}: pixels = 8'b01100110;
            {8'd56, 3'd5}: pixels = 8'b01100110;
            {8'd56, 3'd6}: pixels = 8'b00111100;
            {8'd56, 3'd7}: pixels = 8'b00000000;
            {8'd57, 3'd0}: pixels = 8'b00111100;
            {8'd57, 3'd1}: pixels = 8'b01100110;
            {8'd57, 3'd2}: pixels = 8'b01100110;
            {8'd57, 3'd3}: pixels = 8'b00111110;
            {8'd57, 3'd4}: pixels = 8'b00000110;
            {8'd57, 3'd5}: pixels = 8'b00001100;
            {8'd57, 3'd6}: pixels = 8'b00111000;
            {8'd57, 3'd7}: pixels = 8'b00000000;
            default: pixels = 8'b00000000;
        endcase
    end

endmodule